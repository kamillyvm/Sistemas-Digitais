library verilog;
use verilog.vl_types.all;
entity questao1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        s               : out    vl_logic
    );
end questao1;
