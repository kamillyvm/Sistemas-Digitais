library verilog;
use verilog.vl_types.all;
entity questao2 is
    port(
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        a3              : in     vl_logic;
        s               : out    vl_logic
    );
end questao2;
