library verilog;
use verilog.vl_types.all;
entity questao1_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end questao1_vlg_check_tst;
