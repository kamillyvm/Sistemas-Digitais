library verilog;
use verilog.vl_types.all;
entity questao2_vlg_vec_tst is
end questao2_vlg_vec_tst;
