library verilog;
use verilog.vl_types.all;
entity questao2_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end questao2_vlg_check_tst;
