library verilog;
use verilog.vl_types.all;
entity questao3 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        s1              : out    vl_logic;
        s2              : out    vl_logic
    );
end questao3;
