library verilog;
use verilog.vl_types.all;
entity questao3_vlg_vec_tst is
end questao3_vlg_vec_tst;
