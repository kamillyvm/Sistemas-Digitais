library verilog;
use verilog.vl_types.all;
entity questao1_vlg_vec_tst is
end questao1_vlg_vec_tst;
